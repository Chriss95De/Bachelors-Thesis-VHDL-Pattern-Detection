

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all; 
library altera_mf;
use altera_mf.altera_mf_components.all;

entity WhiteBalance is
port (	

	en				: in std_logic;
	
	amp			: in unsigned(4 downto 0);	
	x_l1			: in unsigned(23 downto 0);
	x_l2			: in unsigned(23 downto 0);
	x_l3			: in unsigned(23 downto 0);
	y_l1			: out unsigned(23 downto 0);
	y_l2			: out unsigned(23 downto 0);
	y_l3			: out unsigned(23 downto 0)
	 
	); 
end entity WhiteBalance;
	
	
architecture a of WhiteBalance is	

	type t_lookuptable is array (0 to 255) of unsigned(7 downto 0);
	
	-- 2
	constant amp_00 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(158,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(166,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(174,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(179,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(184,8),to_unsigned(186,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(191,8),to_unsigned(193,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(198,8),to_unsigned(200,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(205,8),to_unsigned(207,8),to_unsigned(209,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(214,8),to_unsigned(216,8),to_unsigned(218,8),to_unsigned(220,8),to_unsigned(222,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(227,8),to_unsigned(229,8),to_unsigned(231,8),to_unsigned(233,8),to_unsigned(235,8),to_unsigned(237,8),to_unsigned(239,8),to_unsigned(241,8),to_unsigned(243,8),to_unsigned(245,8),to_unsigned(247,8),to_unsigned(249,8),to_unsigned(251,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.9
	constant amp_01 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(168,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(179,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(184,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(192,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(197,8),to_unsigned(199,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(204,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(209,8),to_unsigned(211,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(216,8),to_unsigned(218,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(223,8),to_unsigned(225,8),to_unsigned(227,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(232,8),to_unsigned(234,8),to_unsigned(236,8),to_unsigned(238,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(243,8),to_unsigned(245,8),to_unsigned(247,8),to_unsigned(249,8),to_unsigned(251,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.8
	constant amp_02 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(187,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(195,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(203,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(208,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(213,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(218,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(223,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(228,8),to_unsigned(230,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(235,8),to_unsigned(237,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(242,8),to_unsigned(244,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(249,8),to_unsigned(251,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.7
	constant amp_03 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(201,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(215,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(223,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(228,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(236,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(241,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(246,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(251,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.6
	constant amp_04 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(234,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(245,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.5
	constant amp_05 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.4
	constant amp_06 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.3
	constant amp_07 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.2
	constant amp_08 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1.1
	constant amp_09 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(0,8),to_unsigned(1,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(255,8)
	);
	-- 1
	constant amp_10 : t_lookuptable := (	
	to_unsigned(0,8),to_unsigned(1,8),to_unsigned(2,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(23,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.1
	constant amp_11 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(1,8),to_unsigned(3,8),to_unsigned(4,8),to_unsigned(5,8),to_unsigned(7,8),to_unsigned(8,8),to_unsigned(9,8),to_unsigned(10,8),to_unsigned(12,8),to_unsigned(13,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(20,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(43,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.2
	constant amp_12 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(2,8),to_unsigned(4,8),to_unsigned(6,8),to_unsigned(7,8),to_unsigned(9,8),to_unsigned(11,8),to_unsigned(12,8),to_unsigned(14,8),to_unsigned(15,8),to_unsigned(17,8),to_unsigned(18,8),to_unsigned(19,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(26,8),to_unsigned(27,8),to_unsigned(29,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.3
	constant amp_13 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(3,8),to_unsigned(6,8),to_unsigned(8,8),to_unsigned(10,8),to_unsigned(12,8),to_unsigned(14,8),to_unsigned(16,8),to_unsigned(17,8),to_unsigned(19,8),to_unsigned(21,8),to_unsigned(22,8),to_unsigned(24,8),to_unsigned(25,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(30,8),to_unsigned(31,8),to_unsigned(33,8),to_unsigned(34,8),to_unsigned(35,8),to_unsigned(37,8),to_unsigned(38,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(47,8),to_unsigned(49,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(64,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.4
	constant amp_14 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(4,8),to_unsigned(7,8),to_unsigned(10,8),to_unsigned(13,8),to_unsigned(15,8),to_unsigned(17,8),to_unsigned(19,8),to_unsigned(21,8),to_unsigned(23,8),to_unsigned(25,8),to_unsigned(27,8),to_unsigned(28,8),to_unsigned(30,8),to_unsigned(32,8),to_unsigned(33,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(38,8),to_unsigned(39,8),to_unsigned(41,8),to_unsigned(42,8),to_unsigned(44,8),to_unsigned(45,8),to_unsigned(47,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(53,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(57,8),to_unsigned(59,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.5
	constant amp_15 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(6,8),to_unsigned(10,8),to_unsigned(13,8),to_unsigned(15,8),to_unsigned(18,8),to_unsigned(20,8),to_unsigned(23,8),to_unsigned(25,8),to_unsigned(27,8),to_unsigned(29,8),to_unsigned(31,8),to_unsigned(33,8),to_unsigned(35,8),to_unsigned(36,8),to_unsigned(38,8),to_unsigned(40,8),to_unsigned(41,8),to_unsigned(43,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(48,8),to_unsigned(49,8),to_unsigned(51,8),to_unsigned(52,8),to_unsigned(54,8),to_unsigned(55,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(63,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(67,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(74,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.6
	constant amp_16 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(7,8),to_unsigned(12,8),to_unsigned(15,8),to_unsigned(18,8),to_unsigned(21,8),to_unsigned(24,8),to_unsigned(26,8),to_unsigned(29,8),to_unsigned(31,8),to_unsigned(33,8),to_unsigned(35,8),to_unsigned(37,8),to_unsigned(39,8),to_unsigned(41,8),to_unsigned(43,8),to_unsigned(45,8),to_unsigned(46,8),to_unsigned(48,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(53,8),to_unsigned(55,8),to_unsigned(56,8),to_unsigned(58,8),to_unsigned(59,8),to_unsigned(61,8),to_unsigned(62,8),to_unsigned(64,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(71,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(78,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(83,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.7
	constant amp_17 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(9,8),to_unsigned(14,8),to_unsigned(18,8),to_unsigned(22,8),to_unsigned(25,8),to_unsigned(28,8),to_unsigned(30,8),to_unsigned(33,8),to_unsigned(35,8),to_unsigned(37,8),to_unsigned(40,8),to_unsigned(42,8),to_unsigned(44,8),to_unsigned(46,8),to_unsigned(48,8),to_unsigned(50,8),to_unsigned(51,8),to_unsigned(53,8),to_unsigned(55,8),to_unsigned(57,8),to_unsigned(58,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(63,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(68,8),to_unsigned(69,8),to_unsigned(70,8),to_unsigned(72,8),to_unsigned(73,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.8
	constant amp_18 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(11,8),to_unsigned(17,8),to_unsigned(21,8),to_unsigned(25,8),to_unsigned(28,8),to_unsigned(31,8),to_unsigned(34,8),to_unsigned(37,8),to_unsigned(39,8),to_unsigned(42,8),to_unsigned(44,8),to_unsigned(46,8),to_unsigned(48,8),to_unsigned(50,8),to_unsigned(52,8),to_unsigned(54,8),to_unsigned(56,8),to_unsigned(58,8),to_unsigned(60,8),to_unsigned(61,8),to_unsigned(63,8),to_unsigned(65,8),to_unsigned(67,8),to_unsigned(68,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(76,8),to_unsigned(77,8),to_unsigned(79,8),to_unsigned(80,8),to_unsigned(81,8),to_unsigned(83,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(101,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(106,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/1.9
	constant amp_19 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(13,8),to_unsigned(19,8),to_unsigned(24,8),to_unsigned(28,8),to_unsigned(32,8),to_unsigned(35,8),to_unsigned(38,8),to_unsigned(41,8),to_unsigned(43,8),to_unsigned(46,8),to_unsigned(48,8),to_unsigned(51,8),to_unsigned(53,8),to_unsigned(55,8),to_unsigned(57,8),to_unsigned(59,8),to_unsigned(61,8),to_unsigned(63,8),to_unsigned(65,8),to_unsigned(66,8),to_unsigned(68,8),to_unsigned(70,8),to_unsigned(71,8),to_unsigned(73,8),to_unsigned(75,8),to_unsigned(76,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(86,8),to_unsigned(88,8),to_unsigned(89,8),to_unsigned(91,8),to_unsigned(92,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(96,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(101,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(113,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);
	-- 1/2
	constant amp_20 : t_lookuptable := (	
		to_unsigned(0,8),to_unsigned(15,8),to_unsigned(22,8),to_unsigned(27,8),to_unsigned(31,8),to_unsigned(35,8),to_unsigned(39,8),to_unsigned(42,8),to_unsigned(45,8),to_unsigned(47,8),to_unsigned(50,8),to_unsigned(52,8),to_unsigned(55,8),to_unsigned(57,8),to_unsigned(59,8),to_unsigned(61,8),to_unsigned(63,8),to_unsigned(65,8),to_unsigned(67,8),to_unsigned(69,8),to_unsigned(71,8),to_unsigned(73,8),to_unsigned(74,8),to_unsigned(76,8),to_unsigned(78,8),to_unsigned(79,8),to_unsigned(81,8),to_unsigned(82,8),to_unsigned(84,8),to_unsigned(85,8),to_unsigned(87,8),to_unsigned(88,8),to_unsigned(90,8),to_unsigned(91,8),to_unsigned(93,8),to_unsigned(94,8),to_unsigned(95,8),to_unsigned(97,8),to_unsigned(98,8),to_unsigned(99,8),to_unsigned(100,8),to_unsigned(102,8),to_unsigned(103,8),to_unsigned(104,8),to_unsigned(105,8),to_unsigned(107,8),to_unsigned(108,8),to_unsigned(109,8),to_unsigned(110,8),to_unsigned(111,8),to_unsigned(112,8),to_unsigned(114,8),to_unsigned(115,8),to_unsigned(116,8),to_unsigned(117,8),to_unsigned(118,8),to_unsigned(119,8),to_unsigned(120,8),to_unsigned(121,8),to_unsigned(122,8),to_unsigned(123,8),to_unsigned(124,8),to_unsigned(125,8),to_unsigned(126,8),to_unsigned(127,8),to_unsigned(128,8),to_unsigned(129,8),to_unsigned(130,8),to_unsigned(131,8),to_unsigned(132,8),to_unsigned(133,8),to_unsigned(134,8),to_unsigned(135,8),to_unsigned(136,8),to_unsigned(137,8),to_unsigned(138,8),to_unsigned(139,8),to_unsigned(140,8),to_unsigned(141,8),to_unsigned(141,8),to_unsigned(142,8),to_unsigned(143,8),to_unsigned(144,8),to_unsigned(145,8),to_unsigned(146,8),to_unsigned(147,8),to_unsigned(148,8),to_unsigned(148,8),to_unsigned(149,8),to_unsigned(150,8),to_unsigned(151,8),to_unsigned(152,8),to_unsigned(153,8),to_unsigned(153,8),to_unsigned(154,8),to_unsigned(155,8),to_unsigned(156,8),to_unsigned(157,8),to_unsigned(158,8),to_unsigned(158,8),to_unsigned(159,8),to_unsigned(160,8),to_unsigned(161,8),to_unsigned(162,8),to_unsigned(162,8),to_unsigned(163,8),to_unsigned(164,8),to_unsigned(165,8),to_unsigned(165,8),to_unsigned(166,8),to_unsigned(167,8),to_unsigned(168,8),to_unsigned(168,8),to_unsigned(169,8),to_unsigned(170,8),to_unsigned(171,8),to_unsigned(171,8),to_unsigned(172,8),to_unsigned(173,8),to_unsigned(174,8),to_unsigned(174,8),to_unsigned(175,8),to_unsigned(176,8),to_unsigned(177,8),to_unsigned(177,8),to_unsigned(178,8),to_unsigned(179,8),to_unsigned(179,8),to_unsigned(180,8),to_unsigned(181,8),to_unsigned(182,8),to_unsigned(182,8),to_unsigned(183,8),to_unsigned(184,8),to_unsigned(184,8),to_unsigned(185,8),to_unsigned(186,8),to_unsigned(186,8),to_unsigned(187,8),to_unsigned(188,8),to_unsigned(188,8),to_unsigned(189,8),to_unsigned(190,8),to_unsigned(190,8),to_unsigned(191,8),to_unsigned(192,8),to_unsigned(192,8),to_unsigned(193,8),to_unsigned(194,8),to_unsigned(194,8),to_unsigned(195,8),to_unsigned(196,8),to_unsigned(196,8),to_unsigned(197,8),to_unsigned(198,8),to_unsigned(198,8),to_unsigned(199,8),to_unsigned(200,8),to_unsigned(200,8),to_unsigned(201,8),to_unsigned(201,8),to_unsigned(202,8),to_unsigned(203,8),to_unsigned(203,8),to_unsigned(204,8),to_unsigned(205,8),to_unsigned(205,8),to_unsigned(206,8),to_unsigned(206,8),to_unsigned(207,8),to_unsigned(208,8),to_unsigned(208,8),to_unsigned(209,8),to_unsigned(210,8),to_unsigned(210,8),to_unsigned(211,8),to_unsigned(211,8),to_unsigned(212,8),to_unsigned(213,8),to_unsigned(213,8),to_unsigned(214,8),to_unsigned(214,8),to_unsigned(215,8),to_unsigned(216,8),to_unsigned(216,8),to_unsigned(217,8),to_unsigned(217,8),to_unsigned(218,8),to_unsigned(218,8),to_unsigned(219,8),to_unsigned(220,8),to_unsigned(220,8),to_unsigned(221,8),to_unsigned(221,8),to_unsigned(222,8),to_unsigned(222,8),to_unsigned(223,8),to_unsigned(224,8),to_unsigned(224,8),to_unsigned(225,8),to_unsigned(225,8),to_unsigned(226,8),to_unsigned(226,8),to_unsigned(227,8),to_unsigned(228,8),to_unsigned(228,8),to_unsigned(229,8),to_unsigned(229,8),to_unsigned(230,8),to_unsigned(230,8),to_unsigned(231,8),to_unsigned(231,8),to_unsigned(232,8),to_unsigned(233,8),to_unsigned(233,8),to_unsigned(234,8),to_unsigned(234,8),to_unsigned(235,8),to_unsigned(235,8),to_unsigned(236,8),to_unsigned(236,8),to_unsigned(237,8),to_unsigned(237,8),to_unsigned(238,8),to_unsigned(238,8),to_unsigned(239,8),to_unsigned(240,8),to_unsigned(240,8),to_unsigned(241,8),to_unsigned(241,8),to_unsigned(242,8),to_unsigned(242,8),to_unsigned(243,8),to_unsigned(243,8),to_unsigned(244,8),to_unsigned(244,8),to_unsigned(245,8),to_unsigned(245,8),to_unsigned(246,8),to_unsigned(246,8),to_unsigned(247,8),to_unsigned(247,8),to_unsigned(248,8),to_unsigned(248,8),to_unsigned(249,8),to_unsigned(249,8),to_unsigned(250,8),to_unsigned(250,8),to_unsigned(251,8),to_unsigned(251,8),to_unsigned(252,8),to_unsigned(252,8),to_unsigned(253,8),to_unsigned(253,8),to_unsigned(254,8),to_unsigned(255,8)
	);

	-- Get value from lookup table
	function lookup(x : in unsigned(7 downto 0); a : in unsigned(4 downto 0)) return unsigned is
	begin
		if a = 0 then
			return amp_00(to_integer(x));
		elsif a = 1 then
			return amp_01(to_integer(x));
		elsif a = 2 then
			return amp_02(to_integer(x));
		elsif a = 3 then
			return amp_03(to_integer(x));
		elsif a = 4 then
			return amp_04(to_integer(x));
		elsif a = 5 then
			return amp_05(to_integer(x));
		elsif a = 6 then
			return amp_06(to_integer(x));
		elsif a = 7 then
			return amp_07(to_integer(x));
		elsif a = 8 then
			return amp_08(to_integer(x));
		elsif a = 9 then
			return amp_09(to_integer(x));
		elsif a = 10 then
			return amp_10(to_integer(x));
		elsif a = 11 then
			return amp_11(to_integer(x));
		elsif a = 12 then
			return amp_12(to_integer(x));
		elsif a = 13 then
			return amp_13(to_integer(x));
		elsif a = 14 then
			return amp_14(to_integer(x));
		elsif a = 15 then
			return amp_15(to_integer(x));
		elsif a = 16 then
			return amp_16(to_integer(x));
		elsif a = 17 then
			return amp_17(to_integer(x));
		elsif a = 18 then
			return amp_18(to_integer(x));
		elsif a = 19 then
			return amp_19(to_integer(x));
		elsif a = 20 then
			return amp_20(to_integer(x));
		else
			return amp_10(to_integer(x));
		end if;
	end function;
begin
	
process(en, x_l1, x_l2, x_l3, amp)
begin
	if en = '1' then
		y_l1(23 downto 16) <= lookup(x_l1(23 downto 16), amp);
		y_l1(15 downto 8)  <= lookup(x_l1(15 downto 8), amp);
		y_l1(7 downto 0)   <= lookup(x_l1(7 downto 0), amp);
		y_l2(23 downto 16) <= lookup(x_l2(23 downto 16), amp);
		y_l2(15 downto 8)  <= lookup(x_l2(15 downto 8), amp);
		y_l2(7 downto 0)   <= lookup(x_l2(7 downto 0), amp);
		y_l3(23 downto 16) <= lookup(x_l3(23 downto 16), amp);
		y_l3(15 downto 8)  <= lookup(x_l3(15 downto 8), amp);
		y_l3(7 downto 0)   <= lookup(x_l3(7 downto 0), amp);
	else
		y_l1 <= x_l1;
		y_l2 <= x_l2;
		y_l3 <= x_l3;
	end if;
end process;
end architecture a;